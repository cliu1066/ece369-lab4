`timescale 1ns / 1ps

module ALUControl();

endmodule
